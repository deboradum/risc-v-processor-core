`define ALU_AND         4'b0000
`define ALU_OR          4'b0001
`define ALU_ADD         4'b0010
`define ALU_SUBTRACT    4'b0110
`define ALU_SRL         4'b1000
`define ALU_SLL         4'b1001
`define ALU_SRA         4'b1010

`define RTYPE   7'b0110011
`define LWTYPE   7'b0000011
`define ITYPE   7'b0010011
`define SBTYPE  7'b1100011
`define STYPE   7'b0100011
